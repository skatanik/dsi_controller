// top_level_system_tb.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module top_level_system_tb (
	);

	wire    top_level_system_inst_clk_bfm_clk_clk;       // top_level_system_inst_clk_bfm:clk -> [top_level_system_inst:clk_clk, top_level_system_inst_reset_bfm:clk]
	wire    top_level_system_inst_reset_bfm_reset_reset; // top_level_system_inst_reset_bfm:reset -> top_level_system_inst:reset_reset_n

wire [3:0]	dsi_tx_controller_0_dsi_interface_dphy_data_hs_out_p;
wire [3:0]	dsi_tx_controller_0_dsi_interface_dphy_data_hs_out_n;
wire [3:0]	dsi_tx_controller_0_dsi_interface_dphy_data_lp_out_p;
wire [3:0]	dsi_tx_controller_0_dsi_interface_dphy_data_lp_out_n;
wire 	dsi_tx_controller_0_dsi_interface_dphy_clk_hs_out_p;
wire 	dsi_tx_controller_0_dsi_interface_dphy_clk_hs_out_n;
wire 	dsi_tx_controller_0_dsi_interface_dphy_clk_lp_out_p;
wire 	dsi_tx_controller_0_dsi_interface_dphy_clk_lp_out_n;

	top_level_system top_level_system_inst (
		.altpll_0_areset_conduit_export                       (1'b0),                                            //           altpll_0_areset_conduit.export
		.clk_clk                                              (top_level_system_inst_clk_bfm_clk_clk),       //                               clk.clk
		.dsi_tx_controller_0_dsi_interface_dphy_data_hs_out_p (dsi_tx_controller_0_dsi_interface_dphy_data_hs_out_p ),                                            // dsi_tx_controller_0_dsi_interface.dphy_data_hs_out_p
		.dsi_tx_controller_0_dsi_interface_dphy_data_hs_out_n (dsi_tx_controller_0_dsi_interface_dphy_data_hs_out_n ),                                            //                                  .dphy_data_hs_out_n
		.dsi_tx_controller_0_dsi_interface_dphy_data_lp_out_p (dsi_tx_controller_0_dsi_interface_dphy_data_lp_out_p ),                                            //                                  .dphy_data_lp_out_p
		.dsi_tx_controller_0_dsi_interface_dphy_data_lp_out_n (dsi_tx_controller_0_dsi_interface_dphy_data_lp_out_n ),                                            //                                  .dphy_data_lp_out_n
		.dsi_tx_controller_0_dsi_interface_dphy_clk_hs_out_p  (dsi_tx_controller_0_dsi_interface_dphy_clk_hs_out_p  ),                                            //                                  .dphy_clk_hs_out_p
		.dsi_tx_controller_0_dsi_interface_dphy_clk_hs_out_n  (dsi_tx_controller_0_dsi_interface_dphy_clk_hs_out_n  ),                                            //                                  .dphy_clk_hs_out_n
		.dsi_tx_controller_0_dsi_interface_dphy_clk_lp_out_p  (dsi_tx_controller_0_dsi_interface_dphy_clk_lp_out_p  ),                                            //                                  .dphy_clk_lp_out_p
		.dsi_tx_controller_0_dsi_interface_dphy_clk_lp_out_n  (dsi_tx_controller_0_dsi_interface_dphy_clk_lp_out_n  ),                                            //                                  .dphy_clk_lp_out_n
		.reset_reset_n                                        (top_level_system_inst_reset_bfm_reset_reset)  //                             reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) top_level_system_inst_clk_bfm (
		.clk (top_level_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) top_level_system_inst_reset_bfm (
		.reset (top_level_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (top_level_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
