
mig_ddr3 # (
    .C3_P0_MASK_SIZE(4),
    .C3_P0_DATA_PORT_SIZE(32),
    .C3_P1_MASK_SIZE(4),
    .C3_P1_DATA_PORT_SIZE(32),
    .DEBUG_EN(0),
    .C3_MEMCLK_PERIOD(3000),
    .C3_CALIB_SOFT_IP("TRUE"),
    .C3_SIMULATION("FALSE"),
    .C3_RST_ACT_LOW(0),
    .C3_INPUT_CLK_TYPE("SINGLE_ENDED"),
    .C3_MEM_ADDR_ORDER("BANK_ROW_COLUMN"),
    .C3_NUM_DQ_PINS(16),
    .C3_MEM_ADDR_WIDTH(14),
    .C3_MEM_BANKADDR_WIDTH(3),
    .C3_S0_AXI_STRICT_COHERENCY(0),
    .C3_S0_AXI_ENABLE_AP(0),
    .C3_S0_AXI_DATA_WIDTH(32),
    .C3_S0_AXI_SUPPORTS_NARROW_BURST(1),
    .C3_S0_AXI_ADDR_WIDTH(32),
    .C3_S0_AXI_ID_WIDTH(4),
    .C3_S2_AXI_STRICT_COHERENCY(0),
    .C3_S2_AXI_ENABLE_AP(0),
    .C3_S2_AXI_DATA_WIDTH(32),
    .C3_S2_AXI_SUPPORTS_NARROW_BURST(1),
    .C3_S2_AXI_ADDR_WIDTH(32),
    .C3_S2_AXI_ID_WIDTH(4),
    .C3_S3_AXI_STRICT_COHERENCY(0),
    .C3_S3_AXI_ENABLE_AP(0),
    .C3_S3_AXI_DATA_WIDTH(32),
    .C3_S3_AXI_SUPPORTS_NARROW_BURST(1),
    .C3_S3_AXI_ADDR_WIDTH(32),
    .C3_S3_AXI_ID_WIDTH(4)
)
u_mig_ddr3 (

    .c3_sys_clk           (c3_sys_clk),
  .c3_sys_rst_i           (c3_sys_rst_i),

  .mcb3_dram_dq           (mcb3_dram_dq),
  .mcb3_dram_a            (mcb3_dram_a),
  .mcb3_dram_ba           (mcb3_dram_ba),
  .mcb3_dram_ras_n        (mcb3_dram_ras_n),
  .mcb3_dram_cas_n        (mcb3_dram_cas_n),
  .mcb3_dram_we_n         (mcb3_dram_we_n),
  .mcb3_dram_odt          (mcb3_dram_odt),
  .mcb3_dram_cke          (mcb3_dram_cke),
  .mcb3_dram_ck           (mcb3_dram_ck),
  .mcb3_dram_ck_n         (mcb3_dram_ck_n),
  .mcb3_dram_dqs          (mcb3_dram_dqs),
  .mcb3_dram_dqs_n        (mcb3_dram_dqs_n),
  .mcb3_dram_udqs         (mcb3_dram_udqs),    // for X16 parts
  .mcb3_dram_udqs_n       (mcb3_dram_udqs_n),  // for X16 parts
  .mcb3_dram_udm          (mcb3_dram_udm),     // for X16 parts
  .mcb3_dram_dm           (mcb3_dram_dm),
  .mcb3_dram_reset_n      (mcb3_dram_reset_n),
  .c3_clk0		        (c3_clk0),
  .c3_rst0		        (c3_rst0),



  .c3_calib_done    (c3_calib_done),
     .mcb3_rzq               (rzq3),

     .mcb3_zio               (zio3),

    .c3_s0_axi_aclk                         (c3_s0_axi_aclk   ),
    .c3_s0_axi_aresetn                      (c3_s0_axi_aresetn),
    .c3_s0_axi_awid                         (c3_s0_axi_awid   ),
    .c3_s0_axi_awaddr                       (c3_s0_axi_awaddr ),
    .c3_s0_axi_awlen                        (c3_s0_axi_awlen  ),
    .c3_s0_axi_awsize                       (c3_s0_axi_awsize ),
    .c3_s0_axi_awburst                      (c3_s0_axi_awburst),
    .c3_s0_axi_awlock                       (c3_s0_axi_awlock ),
    .c3_s0_axi_awcache                      (c3_s0_axi_awcache),
    .c3_s0_axi_awprot                       (c3_s0_axi_awprot ),
    .c3_s0_axi_awqos                        (c3_s0_axi_awqos  ),
    .c3_s0_axi_awvalid                      (c3_s0_axi_awvalid),
    .c3_s0_axi_awready                      (c3_s0_axi_awready),
    .c3_s0_axi_wdata                        (c3_s0_axi_wdata  ),
    .c3_s0_axi_wstrb                        (c3_s0_axi_wstrb  ),
    .c3_s0_axi_wlast                        (c3_s0_axi_wlast  ),
    .c3_s0_axi_wvalid                       (c3_s0_axi_wvalid ),
    .c3_s0_axi_wready                       (c3_s0_axi_wready ),
    .c3_s0_axi_bid                          (c3_s0_axi_bid    ),
    .c3_s0_axi_wid                          (c3_s0_axi_wid    ),
    .c3_s0_axi_bresp                        (c3_s0_axi_bresp  ),
    .c3_s0_axi_bvalid                       (c3_s0_axi_bvalid ),
    .c3_s0_axi_bready                       (c3_s0_axi_bready ),
    .c3_s0_axi_arid                         (c3_s0_axi_arid   ),
    .c3_s0_axi_araddr                       (c3_s0_axi_araddr ),
    .c3_s0_axi_arlen                        (c3_s0_axi_arlen  ),
    .c3_s0_axi_arsize                       (c3_s0_axi_arsize ),
    .c3_s0_axi_arburst                      (c3_s0_axi_arburst),
    .c3_s0_axi_arlock                       (c3_s0_axi_arlock ),
    .c3_s0_axi_arcache                      (c3_s0_axi_arcache),
    .c3_s0_axi_arprot                       (c3_s0_axi_arprot ),
    .c3_s0_axi_arqos                        (c3_s0_axi_arqos  ),
    .c3_s0_axi_arvalid                      (c3_s0_axi_arvalid),
    .c3_s0_axi_arready                      (c3_s0_axi_arready),
    .c3_s0_axi_rid                          (c3_s0_axi_rid    ),
    .c3_s0_axi_rdata                        (c3_s0_axi_rdata  ),
    .c3_s0_axi_rresp                        (c3_s0_axi_rresp  ),
    .c3_s0_axi_rlast                        (c3_s0_axi_rlast  ),
    .c3_s0_axi_rvalid                       (c3_s0_axi_rvalid ),
    .c3_s0_axi_rready                       (c3_s0_axi_rready ),

    //* Write only Port
    .c3_s2_axi_aclk                         (c3_s2_axi_aclk   ),
    .c3_s2_axi_aresetn                      (c3_s2_axi_aresetn),
    .c3_s2_axi_awid                         (c3_s2_axi_awid   ),
    .c3_s2_axi_awaddr                       (c3_s2_axi_awaddr ),
    .c3_s2_axi_awlen                        (c3_s2_axi_awlen  ),
    .c3_s2_axi_awsize                       (c3_s2_axi_awsize ),
    .c3_s2_axi_awburst                      (c3_s2_axi_awburst),
    .c3_s2_axi_awlock                       (c3_s2_axi_awlock ),
    .c3_s2_axi_awcache                      (c3_s2_axi_awcache),
    .c3_s2_axi_awprot                       (c3_s2_axi_awprot ),
    .c3_s2_axi_awqos                        (c3_s2_axi_awqos  ),
    .c3_s2_axi_awvalid                      (c3_s2_axi_awvalid),
    .c3_s2_axi_awready                      (c3_s2_axi_awready),
    .c3_s2_axi_wdata                        (c3_s2_axi_wdata  ),
    .c3_s2_axi_wstrb                        (c3_s2_axi_wstrb  ),
    .c3_s2_axi_wlast                        (c3_s2_axi_wlast  ),
    .c3_s2_axi_wvalid                       (c3_s2_axi_wvalid ),
    .c3_s2_axi_wready                       (c3_s2_axi_wready ),
    .c3_s2_axi_bid                          (c3_s2_axi_bid    ),
    .c3_s2_axi_wid                          (c3_s2_axi_wid    ),
    .c3_s2_axi_bresp                        (c3_s2_axi_bresp  ),
    .c3_s2_axi_bvalid                       (c3_s2_axi_bvalid ),
    .c3_s2_axi_bready                       (c3_s2_axi_bready ),
    .c3_s2_axi_arid                         (c3_s2_axi_arid   ),
    .c3_s2_axi_araddr                       (c3_s2_axi_araddr ),
    .c3_s2_axi_arlen                        (c3_s2_axi_arlen  ),
    .c3_s2_axi_arsize                       (c3_s2_axi_arsize ),
    .c3_s2_axi_arburst                      (c3_s2_axi_arburst),
    .c3_s2_axi_arlock                       (c3_s2_axi_arlock ),
    .c3_s2_axi_arcache                      (c3_s2_axi_arcache),
    .c3_s2_axi_arprot                       (c3_s2_axi_arprot ),
    .c3_s2_axi_arqos                        (c3_s2_axi_arqos  ),
    .c3_s2_axi_arvalid                      (c3_s2_axi_arvalid),
    .c3_s2_axi_arready                      (c3_s2_axi_arready),
    .c3_s2_axi_rid                          (c3_s2_axi_rid    ),
    .c3_s2_axi_rdata                        (c3_s2_axi_rdata  ),
    .c3_s2_axi_rresp                        (c3_s2_axi_rresp  ),
    .c3_s2_axi_rlast                        (c3_s2_axi_rlast  ),
    .c3_s2_axi_rvalid                       (c3_s2_axi_rvalid ),
    .c3_s2_axi_rready                       (c3_s2_axi_rready ),

    //* Read only Port
    .c3_s3_axi_aclk                         (c3_s3_axi_aclk   ),
    .c3_s3_axi_aresetn                      (c3_s3_axi_aresetn),
    .c3_s3_axi_awid                         (c3_s3_axi_awid   ),
    .c3_s3_axi_awaddr                       (c3_s3_axi_awaddr ),
    .c3_s3_axi_awlen                        (c3_s3_axi_awlen  ),
    .c3_s3_axi_awsize                       (c3_s3_axi_awsize ),
    .c3_s3_axi_awburst                      (c3_s3_axi_awburst),
    .c3_s3_axi_awlock                       (c3_s3_axi_awlock ),
    .c3_s3_axi_awcache                      (c3_s3_axi_awcache),
    .c3_s3_axi_awprot                       (c3_s3_axi_awprot ),
    .c3_s3_axi_awqos                        (c3_s3_axi_awqos  ),
    .c3_s3_axi_awvalid                      (c3_s3_axi_awvalid),
    .c3_s3_axi_awready                      (c3_s3_axi_awready),
    .c3_s3_axi_wdata                        (c3_s3_axi_wdata  ),
    .c3_s3_axi_wstrb                        (c3_s3_axi_wstrb  ),
    .c3_s3_axi_wlast                        (c3_s3_axi_wlast  ),
    .c3_s3_axi_wvalid                       (c3_s3_axi_wvalid ),
    .c3_s3_axi_wready                       (c3_s3_axi_wready ),
    .c3_s3_axi_bid                          (c3_s3_axi_bid    ),
    .c3_s3_axi_wid                          (c3_s3_axi_wid    ),
    .c3_s3_axi_bresp                        (c3_s3_axi_bresp  ),
    .c3_s3_axi_bvalid                       (c3_s3_axi_bvalid ),
    .c3_s3_axi_bready                       (c3_s3_axi_bready ),
    .c3_s3_axi_arid                         (c3_s3_axi_arid   ),
    .c3_s3_axi_araddr                       (c3_s3_axi_araddr ),
    .c3_s3_axi_arlen                        (c3_s3_axi_arlen  ),
    .c3_s3_axi_arsize                       (c3_s3_axi_arsize ),
    .c3_s3_axi_arburst                      (c3_s3_axi_arburst),
    .c3_s3_axi_arlock                       (c3_s3_axi_arlock ),
    .c3_s3_axi_arcache                      (c3_s3_axi_arcache),
    .c3_s3_axi_arprot                       (c3_s3_axi_arprot ),
    .c3_s3_axi_arqos                        (c3_s3_axi_arqos  ),
    .c3_s3_axi_arvalid                      (c3_s3_axi_arvalid),
    .c3_s3_axi_arready                      (c3_s3_axi_arready),
    .c3_s3_axi_rid                          (c3_s3_axi_rid    ),
    .c3_s3_axi_rdata                        (c3_s3_axi_rdata  ),
    .c3_s3_axi_rresp                        (c3_s3_axi_rresp  ),
    .c3_s3_axi_rlast                        (c3_s3_axi_rlast  ),
    .c3_s3_axi_rvalid                       (c3_s3_axi_rvalid ),
    .c3_s3_axi_rready                       (c3_s3_axi_rready )
);