`ifndef PRJ_DEFINES
`define PRJ_DEFINES

`define SIMULATION

`endif